module FM_Module(
	input clk,
	input rst,
	input [11:0] dac_modu_12bit,
	output [63:0]freq
);


